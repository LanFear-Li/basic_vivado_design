module decoder_tb_3_to_8;
    
    reg [2:0] A;
    reg STA, STB, STC;
    wire [7:0] Y;
    
    decoder_3_to_8 test(.A(A), .STA(STA), .STB(STB), .STC(STC), .Y(Y));
    
    initial begin
        
        STA = 1;
        STB = 0;
        STC = 0;
        
        A[0] = 0;
        A[1] = 0;
        A[2] = 0;
        #5;
        
        A[0] = 1;
        A[1] = 0;
        A[2] = 0;
        #5;
        
        A[0] = 0;
        A[1] = 1;
        A[2] = 0;
        #5;
        
        A[0] = 1;
        A[1] = 1;
        A[2] = 0;
        #5;
        
        A[0] = 0;
        A[1] = 0;
        A[2] = 1;
        #5;
        
        A[0] = 1;
        A[1] = 0;
        A[2] = 1;
        #5;
        
        A[0] = 0;
        A[1] = 1;
        A[2] = 1;
        #5;
        
        A[0] = 1;
        A[1] = 1;
        A[2] = 1;
        #5;
    end

endmodule

module decoder_tb_4_to_16();
    reg [3:0] A;
    wire [15:0] Y;
    decoder_4_to_16 test(.A(A), .Y(Y));
    
    initial begin
        A[0] = 0;
        A[1] = 0;
        A[2] = 0;
        A[3] = 0;
        #5;
        
        A[0] = 1;
        A[1] = 0;
        A[2] = 0;
        A[3] = 0;
        #5;
        A[0] = 0;
        A[1] = 1;
        A[2] = 0;
        A[3] = 0;
        #5;
        
        A[0] = 1;
        A[1] = 1;
        A[2] = 0;
        A[3] = 0;
        #5;
        
        A[0] = 0;
        A[1] = 0;
        A[2] = 1;
        A[3] = 0;
        #5;
        
        A[0] = 1;
        A[1] = 0;
        A[2] = 1;
        A[3] = 0;
        #5;
        
        A[0] = 0;
        A[1] = 1;
        A[2] = 1;
        A[3] = 0;
        #5;
        
        A[0] = 1;
        A[1] = 1;
        A[2] = 1;
        A[3] = 0;
        #5;
        
        A[0] = 0;
        A[1] = 0;
        A[2] = 0;
        A[3] = 1;
        #5;
        
        A[0] = 1;
        A[1] = 0;
        A[2] = 0;
        A[3] = 1;
        #5;
        
        A[0] = 0;
        A[1] = 1;
        A[2] = 0;
        A[3] = 1;
        #5;
        
        A[0] = 1;
        A[1] = 1;
        A[2] = 0;
        A[3] = 1;
        #5;
        
        A[0] = 0;
        A[1] = 0;
        A[2] = 1;
        A[3] = 1;
        #5;
        
        A[0] = 1;
        A[1] = 0;
        A[2] = 1;
        A[3] = 1;
        #5;
        
        A[0] = 0;
        A[1] = 1;
        A[2] = 1;
        A[3] = 1;
        #5;
        
        A[0] = 1;
        A[1] = 1;
        A[2] = 1;
        A[3] = 1;
        #5;
    end
endmodule